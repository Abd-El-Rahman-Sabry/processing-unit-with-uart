`include "./../parameters.v"

module system_ctrl(
    input wire i_clk , i_rst, 
);

endmodule 